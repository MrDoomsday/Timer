module timer #(
    parameter FREQUENCY_VALUE = 50_000_000//in Hz
) (
    input logic clk,
    input logic reset_n,

    input 	logic   [1:0]	avmms_address,
	input 	logic			avmms_write,
	input 	logic	[31:0]	avmms_writedata,
    input   logic   [3:0]   avmms_byteenable, 
	input 	logic			avmms_read,
	output 	logic 	[31:0]	avmms_readdata,

    output  logic           coe_interrupt
);

/***************************************************************************************************************************/
/***************************************************************************************************************************/
/******************************************								   *************************************************/
/******************************************								   *************************************************/
/******************************************				Declaration		   *************************************************/
/******************************************								   *************************************************/
/******************************************								   *************************************************/
/***************************************************************************************************************************/
/***************************************************************************************************************************/


logic [63:0] counter, counter_reg;
logic complete;
logic busy;
logic start;
logic stop;




/***************************************************************************************************************************/
/***************************************************************************************************************************/
/******************************************								   *************************************************/
/******************************************								   *************************************************/
/******************************************				Avalon-MM		   *************************************************/
/******************************************								   *************************************************/
/******************************************								   *************************************************/
/***************************************************************************************************************************/
/***************************************************************************************************************************/
//ADDRESS = 0
always_ff @ (posedge clk or negedge reset_n)
    if(!reset_n) {stop, start} <= 2'h0;
    else if(avmms_write && (avmms_address == 2'h0)) begin
        if(avmms_byteenable[0]) {stop, start} <= avmms_writedata[1:0];
    end
    else {stop, start} <= 2'h0;



always_ff @ (posedge clk or negedge reset_n)
    if(!reset_n) counter_reg[31:0] <= 32'h0;
    else if(avmms_write && (avmms_address == 2'h1)) begin
        if(avmms_byteenable[3]) counter_reg[31:24] <= avmms_writedata[31:24];
        if(avmms_byteenable[2]) counter_reg[23:16] <= avmms_writedata[23:16];
        if(avmms_byteenable[1]) counter_reg[15:8] <= avmms_writedata[15:8];
        if(avmms_byteenable[0]) counter_reg[7:0] <= avmms_writedata[7:0];
    end

always_ff @ (posedge clk or negedge reset_n)
    if(!reset_n) counter_reg[63:32] <= 32'h0;
    else if(avmms_write && (avmms_address == 2'h2)) begin
        if(avmms_byteenable[3]) counter_reg[63:56] <= avmms_writedata[31:24];
        if(avmms_byteenable[2]) counter_reg[55:48] <= avmms_writedata[23:16];
        if(avmms_byteenable[1]) counter_reg[47:40] <= avmms_writedata[15:8];
        if(avmms_byteenable[0]) counter_reg[39:32] <= avmms_writedata[7:0];
    end

always_ff @ (posedge clk) begin
    case(avmms_address)
        2'h0: avmms_readdata <= {28'h0, complete, busy, stop, start};
        2'h1: avmms_readdata <= counter_reg[31:0];
        2'h2: avmms_readdata <= counter_reg[63:32];
        2'h3: avmms_readdata <= 32'h0;
        default: avmms_readdata <= 32'h0;
    endcase
end

/***************************************************************************************************************************/
/***************************************************************************************************************************/
/******************************************								   *************************************************/
/******************************************								   *************************************************/
/******************************************				Logic   		   *************************************************/
/******************************************								   *************************************************/
/******************************************								   *************************************************/
/***************************************************************************************************************************/
/***************************************************************************************************************************/
always_ff @ (posedge clk or negedge reset_n)
    if(!reset_n) counter <= 64'h0;
    else if(start && (counter_reg > 64'h0)) counter <= counter_reg;
    else if(stop) counter <= 64'h0;
    else if(counter > 64'h0) counter <= counter - 64'h1;

always_ff @ (posedge clk or negedge reset_n)
    if(!reset_n) complete <= 1'b0;
    else if(counter == 64'h1) complete <= 1'b1;
    else if(avmms_write && (avmms_address == 2'h0)) complete <= 1'b0;

always_ff @ (posedge clk or negedge reset_n)
    if(!reset_n) busy <= 1'b0;
    else if(start && (counter_reg > 64'h0)) busy <= 1'b1;
    else if(stop && (counter == 64'h1)) busy <= 1'b0;

assign coe_interrupt = complete;

endmodule